module cubase2_dongle (
	input clk,
	input reset, // POR actually
	input uds_n,
	input [8:1] A,
	output reg [15:8] D
);

reg uds_nD;
always @(posedge clk) begin
	uds_nD <= uds_n;
	if (reset) begin
		D <= 0;
	end
	else
	if (uds_n & !uds_nD) begin
		D[15] <= !( (A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1])
		          | (         D[14] &  D[12]               &  D[10]                    & A[1] )
		          | (                D[13]               & !D[10]             & A[4] )
		          | ( !D[15] & !D[14] & !D[13] & !D[12] & !D[11] &  D[10] & !D[9]       & A[4] )
		          | (        !D[14]                      & !D[10]                    & A[1])
		          | (  D[15]                             & !D[10]             & A[4]  )
		          | (                      !D[12]        & !D[10]                    & A[1])
		          | (  !D[8] & A[5]));

		D[14] <= !((A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1] )
		          | ( !D[15] & !D[14] & !D[13] & !D[12] & !D[11] & !D[10] & !D[9] &  D[8] & A[4])
		          | (         D[14]        &  D[12]        &  D[10]       &  D[8]        & A[1] )
		          | (                                    !D[10]       & !D[8]        & A[1] )
		          | (                      !D[12]                     & !D[8]        & A[1] )
		          | (  D[15]                                          & !D[8] & A[4])
		          | (        !D[14]                                   & !D[8]        & A[1] )
		          | ( !D[15] & A[5]));

		D[13] <= !((A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1] )
		          | (  D[15] &  D[14] &  D[13] &  D[12] &  D[11] &  D[10]       &  D[8]        & A[1] )
		          | ( !D[15]        & !D[13]        &  D[11]                    & A[4] )
		          | (                D[13]        & !D[11]                    & A[4] )
		          | (                      !D[12] & !D[11]                           & A[1]  )
		          | (  D[15]                      & !D[11]                    & A[4] )
		          | (        !D[14]               & !D[11]                           & A[1]  )
		          | ( !D[9] & A[5]));

		D[12] <= !((A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1])
		          | (  D[15] &  D[14] &  D[13] &  D[12]        &  D[10]       &  D[8]        & A[1] )
		          | (               !D[13]               & !D[10]                    & A[1]  )
		          | ( !D[15]        &  D[13]                                  & A[4]  )
		          | (               !D[13] & !D[12]                                  & A[1]  )
		          | (  D[15]        & !D[13]                                  & A[4] )
		          | (        !D[14] & !D[13]                                         & A[1] )
		          | ( !D[11] & A[5]));

		D[11] <= !((A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1])
		          | (  D[15] &  D[14]        &  D[12]        &  D[10]       &  D[8]        & A[1] )
		          | ( !D[15]                                          & !D[8]        & A[1] )
		          | ( !D[15]                             & !D[10]                    & A[1] )
		          | ( !D[15]               & !D[12]                                  & A[1] )
		          | ( !D[15] & !D[14]                                                & A[1] )
		          | (  D[15]                                                & A[4] )
		          | ( !D[13] & A[5]));

		D[10] <= !((A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1] )
		          | (  D[15] &  D[14] &  D[13] &  D[12] &  D[11] &  D[10] &  D[9] &  D[8]        & A[1] )
		          | ( !D[15]        & !D[13]        & !D[11]        &  D[9]       & A[4] )
		          | (                              D[11]        & !D[9]       & A[4] )
		          | (                D[13]                      & !D[9]       & A[4] )
		          | (  D[15]                                    & !D[9]       & A[4] )
		          | (        !D[14] & !D[9]                                          & A[1] )
		          | ( !D[14] & A[5]));

		D[9]  <= !((A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1] )
		          | ( !D[15] &  D[14] & !D[13]         & !D[11]       & !D[9]       & A[4] )
		          | (        !D[14]                             &  D[9]       & A[4] )
		          | (        !D[14]                &  D[11]                   & A[4] )
		          | (        !D[14] &  D[13]                                  & A[4] )
		          | (  D[15] & !D[14]                                         & A[4] )
		          | (         D[14]                                                & A[1] )
		          | ( !D[12] & A[5]));

		D[8] <= !((A[8] & A[7] & !A[6] & A[5] & A[4] & !A[3] & !A[2] & !A[1] )
		          | ( !D[15] & !D[14] & !D[13] &  D[12] & !D[11]        & !D[9]       & A[4] )
		          | (         D[14]        &  D[12]                                  & A[1] )
		          | (                      !D[12] &  D[11]                    & A[4] )
		          | (                D[13] & !D[12]                           & A[4] )
		          | (  D[15]               & !D[12]                           & A[4] )
		          | (       !D[14]         & !D[12]                                  & A[1] )
		          | ( !D[10] & A[5]	));
	end

end

endmodule
