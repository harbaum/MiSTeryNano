module font_8x8_fnt (
  input clk,
  input [10:0] addr,
  output reg [7:0] dout
);

always @( posedge clk) begin
  case (addr)
    11'h000: dout = 8'h00;
    11'h001: dout = 8'h00;
    11'h002: dout = 8'h00;
    11'h003: dout = 8'h00;
    11'h004: dout = 8'h00;
    11'h005: dout = 8'h00;
    11'h006: dout = 8'h00;
    11'h007: dout = 8'h00;
    11'h008: dout = 8'h7e;
    11'h009: dout = 8'h81;
    11'h00a: dout = 8'ha5;
    11'h00b: dout = 8'h81;
    11'h00c: dout = 8'hbd;
    11'h00d: dout = 8'h99;
    11'h00e: dout = 8'h81;
    11'h00f: dout = 8'h7e;
    11'h010: dout = 8'h7e;
    11'h011: dout = 8'hff;
    11'h012: dout = 8'hdb;
    11'h013: dout = 8'hff;
    11'h014: dout = 8'hff;
    11'h015: dout = 8'hc3;
    11'h016: dout = 8'he7;
    11'h017: dout = 8'h7e;
    11'h018: dout = 8'h00;
    11'h019: dout = 8'hee;
    11'h01a: dout = 8'hfe;
    11'h01b: dout = 8'hfe;
    11'h01c: dout = 8'h7c;
    11'h01d: dout = 8'h38;
    11'h01e: dout = 8'h10;
    11'h01f: dout = 8'h00;
    11'h020: dout = 8'h10;
    11'h021: dout = 8'h38;
    11'h022: dout = 8'h7c;
    11'h023: dout = 8'hfe;
    11'h024: dout = 8'h7c;
    11'h025: dout = 8'h38;
    11'h026: dout = 8'h10;
    11'h027: dout = 8'h00;
    11'h028: dout = 8'h18;
    11'h029: dout = 8'h3c;
    11'h02a: dout = 8'h18;
    11'h02b: dout = 8'hff;
    11'h02c: dout = 8'hff;
    11'h02d: dout = 8'h4a;
    11'h02e: dout = 8'h18;
    11'h02f: dout = 8'h00;
    11'h030: dout = 8'h10;
    11'h031: dout = 8'h38;
    11'h032: dout = 8'h7c;
    11'h033: dout = 8'hfe;
    11'h034: dout = 8'hfe;
    11'h035: dout = 8'h92;
    11'h036: dout = 8'h38;
    11'h037: dout = 8'h00;
    11'h038: dout = 8'h00;
    11'h039: dout = 8'h00;
    11'h03a: dout = 8'h18;
    11'h03b: dout = 8'h3c;
    11'h03c: dout = 8'h18;
    11'h03d: dout = 8'h00;
    11'h03e: dout = 8'h00;
    11'h03f: dout = 8'h00;
    11'h040: dout = 8'hff;
    11'h041: dout = 8'hff;
    11'h042: dout = 8'he7;
    11'h043: dout = 8'hc3;
    11'h044: dout = 8'he7;
    11'h045: dout = 8'hff;
    11'h046: dout = 8'hff;
    11'h047: dout = 8'hff;
    11'h048: dout = 8'h00;
    11'h049: dout = 8'h3c;
    11'h04a: dout = 8'h42;
    11'h04b: dout = 8'h81;
    11'h04c: dout = 8'h81;
    11'h04d: dout = 8'h42;
    11'h04e: dout = 8'h3c;
    11'h04f: dout = 8'h00;
    11'h050: dout = 8'hff;
    11'h051: dout = 8'hc3;
    11'h052: dout = 8'hbd;
    11'h053: dout = 8'h7e;
    11'h054: dout = 8'h7e;
    11'h055: dout = 8'hbd;
    11'h056: dout = 8'hc3;
    11'h057: dout = 8'hff;
    11'h058: dout = 8'h1f;
    11'h059: dout = 8'h07;
    11'h05a: dout = 8'h0d;
    11'h05b: dout = 8'h7c;
    11'h05c: dout = 8'hc6;
    11'h05d: dout = 8'hc6;
    11'h05e: dout = 8'h7c;
    11'h05f: dout = 8'h00;
    11'h060: dout = 8'h00;
    11'h061: dout = 8'h7e;
    11'h062: dout = 8'hc3;
    11'h063: dout = 8'hc3;
    11'h064: dout = 8'h7e;
    11'h065: dout = 8'h18;
    11'h066: dout = 8'h7e;
    11'h067: dout = 8'h18;
    11'h068: dout = 8'h04;
    11'h069: dout = 8'h06;
    11'h06a: dout = 8'h07;
    11'h06b: dout = 8'h04;
    11'h06c: dout = 8'h04;
    11'h06d: dout = 8'hfc;
    11'h06e: dout = 8'hf8;
    11'h06f: dout = 8'h00;
    11'h070: dout = 8'h0c;
    11'h071: dout = 8'h0a;
    11'h072: dout = 8'h0d;
    11'h073: dout = 8'h0b;
    11'h074: dout = 8'hf9;
    11'h075: dout = 8'hf1;
    11'h076: dout = 8'h0f;
    11'h077: dout = 8'h0f;
    11'h078: dout = 8'h81;
    11'h079: dout = 8'h43;
    11'h07a: dout = 8'h3d;
    11'h07b: dout = 8'h27;
    11'h07c: dout = 8'h25;
    11'h07d: dout = 8'h3f;
    11'h07e: dout = 8'h57;
    11'h07f: dout = 8'hff;
    11'h080: dout = 8'h00;
    11'h081: dout = 8'h00;
    11'h082: dout = 8'h60;
    11'h083: dout = 8'h78;
    11'h084: dout = 8'h7e;
    11'h085: dout = 8'h78;
    11'h086: dout = 8'h60;
    11'h087: dout = 8'h00;
    11'h088: dout = 8'h00;
    11'h089: dout = 8'h00;
    11'h08a: dout = 8'h06;
    11'h08b: dout = 8'h1e;
    11'h08c: dout = 8'h7e;
    11'h08d: dout = 8'h1e;
    11'h08e: dout = 8'h06;
    11'h08f: dout = 8'h00;
    11'h090: dout = 8'h18;
    11'h091: dout = 8'h7e;
    11'h092: dout = 8'h18;
    11'h093: dout = 8'h18;
    11'h094: dout = 8'h18;
    11'h095: dout = 8'h18;
    11'h096: dout = 8'h7e;
    11'h097: dout = 8'h18;
    11'h098: dout = 8'h66;
    11'h099: dout = 8'h66;
    11'h09a: dout = 8'h66;
    11'h09b: dout = 8'h66;
    11'h09c: dout = 8'h66;
    11'h09d: dout = 8'h00;
    11'h09e: dout = 8'h66;
    11'h09f: dout = 8'h00;
    11'h0a0: dout = 8'hff;
    11'h0a1: dout = 8'hb6;
    11'h0a2: dout = 8'h76;
    11'h0a3: dout = 8'h36;
    11'h0a4: dout = 8'h36;
    11'h0a5: dout = 8'h36;
    11'h0a6: dout = 8'h36;
    11'h0a7: dout = 8'h00;
    11'h0a8: dout = 8'h7e;
    11'h0a9: dout = 8'h81;
    11'h0aa: dout = 8'h7c;
    11'h0ab: dout = 8'h42;
    11'h0ac: dout = 8'h42;
    11'h0ad: dout = 8'h3e;
    11'h0ae: dout = 8'h81;
    11'h0af: dout = 8'h7e;
    11'h0b0: dout = 8'h00;
    11'h0b1: dout = 8'h00;
    11'h0b2: dout = 8'h00;
    11'h0b3: dout = 8'h7e;
    11'h0b4: dout = 8'h7e;
    11'h0b5: dout = 8'h00;
    11'h0b6: dout = 8'h00;
    11'h0b7: dout = 8'h00;
    11'h0b8: dout = 8'h18;
    11'h0b9: dout = 8'h7e;
    11'h0ba: dout = 8'h18;
    11'h0bb: dout = 8'h18;
    11'h0bc: dout = 8'h7e;
    11'h0bd: dout = 8'h18;
    11'h0be: dout = 8'h00;
    11'h0bf: dout = 8'hff;
    11'h0c0: dout = 8'h18;
    11'h0c1: dout = 8'h7e;
    11'h0c2: dout = 8'h18;
    11'h0c3: dout = 8'h18;
    11'h0c4: dout = 8'h18;
    11'h0c5: dout = 8'h18;
    11'h0c6: dout = 8'h18;
    11'h0c7: dout = 8'h00;
    11'h0c8: dout = 8'h18;
    11'h0c9: dout = 8'h18;
    11'h0ca: dout = 8'h18;
    11'h0cb: dout = 8'h18;
    11'h0cc: dout = 8'h18;
    11'h0cd: dout = 8'h7e;
    11'h0ce: dout = 8'h18;
    11'h0cf: dout = 8'h00;
    11'h0d0: dout = 8'h00;
    11'h0d1: dout = 8'h04;
    11'h0d2: dout = 8'h06;
    11'h0d3: dout = 8'hff;
    11'h0d4: dout = 8'h06;
    11'h0d5: dout = 8'h04;
    11'h0d6: dout = 8'h00;
    11'h0d7: dout = 8'h00;
    11'h0d8: dout = 8'h00;
    11'h0d9: dout = 8'h20;
    11'h0da: dout = 8'h60;
    11'h0db: dout = 8'hff;
    11'h0dc: dout = 8'h60;
    11'h0dd: dout = 8'h20;
    11'h0de: dout = 8'h00;
    11'h0df: dout = 8'h00;
    11'h0e0: dout = 8'h00;
    11'h0e1: dout = 8'h00;
    11'h0e2: dout = 8'h00;
    11'h0e3: dout = 8'hc0;
    11'h0e4: dout = 8'hc0;
    11'h0e5: dout = 8'hc0;
    11'h0e6: dout = 8'hff;
    11'h0e7: dout = 8'h00;
    11'h0e8: dout = 8'h00;
    11'h0e9: dout = 8'h24;
    11'h0ea: dout = 8'h66;
    11'h0eb: dout = 8'hff;
    11'h0ec: dout = 8'h66;
    11'h0ed: dout = 8'h24;
    11'h0ee: dout = 8'h00;
    11'h0ef: dout = 8'h00;
    11'h0f0: dout = 8'h00;
    11'h0f1: dout = 8'h00;
    11'h0f2: dout = 8'h10;
    11'h0f3: dout = 8'h38;
    11'h0f4: dout = 8'h7c;
    11'h0f5: dout = 8'hfe;
    11'h0f6: dout = 8'h00;
    11'h0f7: dout = 8'h00;
    11'h0f8: dout = 8'h00;
    11'h0f9: dout = 8'h00;
    11'h0fa: dout = 8'h00;
    11'h0fb: dout = 8'hfe;
    11'h0fc: dout = 8'h7c;
    11'h0fd: dout = 8'h38;
    11'h0fe: dout = 8'h10;
    11'h0ff: dout = 8'h00;
    11'h100: dout = 8'h00;
    11'h101: dout = 8'h00;
    11'h102: dout = 8'h00;
    11'h103: dout = 8'h00;
    11'h104: dout = 8'h00;
    11'h105: dout = 8'h00;
    11'h106: dout = 8'h00;
    11'h107: dout = 8'h00;
    11'h108: dout = 8'h30;
    11'h109: dout = 8'h78;
    11'h10a: dout = 8'h78;
    11'h10b: dout = 8'h78;
    11'h10c: dout = 8'h30;
    11'h10d: dout = 8'h00;
    11'h10e: dout = 8'h30;
    11'h10f: dout = 8'h00;
    11'h110: dout = 8'hcc;
    11'h111: dout = 8'h66;
    11'h112: dout = 8'h33;
    11'h113: dout = 8'h00;
    11'h114: dout = 8'h00;
    11'h115: dout = 8'h00;
    11'h116: dout = 8'h00;
    11'h117: dout = 8'h00;
    11'h118: dout = 8'h00;
    11'h119: dout = 8'h36;
    11'h11a: dout = 8'h7f;
    11'h11b: dout = 8'h36;
    11'h11c: dout = 8'h36;
    11'h11d: dout = 8'h7f;
    11'h11e: dout = 8'h36;
    11'h11f: dout = 8'h00;
    11'h120: dout = 8'h7c;
    11'h121: dout = 8'hd6;
    11'h122: dout = 8'hd0;
    11'h123: dout = 8'h7c;
    11'h124: dout = 8'h16;
    11'h125: dout = 8'hd6;
    11'h126: dout = 8'h7c;
    11'h127: dout = 8'h10;
    11'h128: dout = 8'he3;
    11'h129: dout = 8'ha6;
    11'h12a: dout = 8'hec;
    11'h12b: dout = 8'h18;
    11'h12c: dout = 8'h37;
    11'h12d: dout = 8'h65;
    11'h12e: dout = 8'hc7;
    11'h12f: dout = 8'h00;
    11'h130: dout = 8'h38;
    11'h131: dout = 8'h4c;
    11'h132: dout = 8'h38;
    11'h133: dout = 8'h45;
    11'h134: dout = 8'hc6;
    11'h135: dout = 8'hce;
    11'h136: dout = 8'h7a;
    11'h137: dout = 8'h01;
    11'h138: dout = 8'h06;
    11'h139: dout = 8'h0c;
    11'h13a: dout = 8'h18;
    11'h13b: dout = 8'h00;
    11'h13c: dout = 8'h00;
    11'h13d: dout = 8'h00;
    11'h13e: dout = 8'h00;
    11'h13f: dout = 8'h00;
    11'h140: dout = 8'h0c;
    11'h141: dout = 8'h18;
    11'h142: dout = 8'h18;
    11'h143: dout = 8'h18;
    11'h144: dout = 8'h18;
    11'h145: dout = 8'h18;
    11'h146: dout = 8'h18;
    11'h147: dout = 8'h0c;
    11'h148: dout = 8'h60;
    11'h149: dout = 8'h30;
    11'h14a: dout = 8'h30;
    11'h14b: dout = 8'h30;
    11'h14c: dout = 8'h30;
    11'h14d: dout = 8'h30;
    11'h14e: dout = 8'h30;
    11'h14f: dout = 8'h60;
    11'h150: dout = 8'h10;
    11'h151: dout = 8'h54;
    11'h152: dout = 8'h38;
    11'h153: dout = 8'hfe;
    11'h154: dout = 8'h38;
    11'h155: dout = 8'h54;
    11'h156: dout = 8'h10;
    11'h157: dout = 8'h00;
    11'h158: dout = 8'h00;
    11'h159: dout = 8'h18;
    11'h15a: dout = 8'h18;
    11'h15b: dout = 8'h7e;
    11'h15c: dout = 8'h18;
    11'h15d: dout = 8'h18;
    11'h15e: dout = 8'h00;
    11'h15f: dout = 8'h00;
    11'h160: dout = 8'h00;
    11'h161: dout = 8'h00;
    11'h162: dout = 8'h00;
    11'h163: dout = 8'h00;
    11'h164: dout = 8'h00;
    11'h165: dout = 8'h00;
    11'h166: dout = 8'h18;
    11'h167: dout = 8'h30;
    11'h168: dout = 8'h00;
    11'h169: dout = 8'h00;
    11'h16a: dout = 8'h00;
    11'h16b: dout = 8'h7e;
    11'h16c: dout = 8'h00;
    11'h16d: dout = 8'h00;
    11'h16e: dout = 8'h00;
    11'h16f: dout = 8'h00;
    11'h170: dout = 8'h00;
    11'h171: dout = 8'h00;
    11'h172: dout = 8'h00;
    11'h173: dout = 8'h00;
    11'h174: dout = 8'h00;
    11'h175: dout = 8'h00;
    11'h176: dout = 8'h30;
    11'h177: dout = 8'h00;
    11'h178: dout = 8'h00;
    11'h179: dout = 8'h03;
    11'h17a: dout = 8'h06;
    11'h17b: dout = 8'h0c;
    11'h17c: dout = 8'h18;
    11'h17d: dout = 8'h30;
    11'h17e: dout = 8'h60;
    11'h17f: dout = 8'h00;
    11'h180: dout = 8'h7c;
    11'h181: dout = 8'hce;
    11'h182: dout = 8'hde;
    11'h183: dout = 8'hfe;
    11'h184: dout = 8'hee;
    11'h185: dout = 8'hce;
    11'h186: dout = 8'h7c;
    11'h187: dout = 8'h00;
    11'h188: dout = 8'h1c;
    11'h189: dout = 8'h3c;
    11'h18a: dout = 8'h1c;
    11'h18b: dout = 8'h1c;
    11'h18c: dout = 8'h1c;
    11'h18d: dout = 8'h1c;
    11'h18e: dout = 8'h1c;
    11'h18f: dout = 8'h00;
    11'h190: dout = 8'h7c;
    11'h191: dout = 8'hce;
    11'h192: dout = 8'h0e;
    11'h193: dout = 8'h1c;
    11'h194: dout = 8'h38;
    11'h195: dout = 8'h70;
    11'h196: dout = 8'hfe;
    11'h197: dout = 8'h00;
    11'h198: dout = 8'h7c;
    11'h199: dout = 8'hce;
    11'h19a: dout = 8'h0e;
    11'h19b: dout = 8'h3c;
    11'h19c: dout = 8'h0e;
    11'h19d: dout = 8'hce;
    11'h19e: dout = 8'h7c;
    11'h19f: dout = 8'h00;
    11'h1a0: dout = 8'hce;
    11'h1a1: dout = 8'hce;
    11'h1a2: dout = 8'hce;
    11'h1a3: dout = 8'hce;
    11'h1a4: dout = 8'hfe;
    11'h1a5: dout = 8'h0e;
    11'h1a6: dout = 8'h0e;
    11'h1a7: dout = 8'h00;
    11'h1a8: dout = 8'hfe;
    11'h1a9: dout = 8'he0;
    11'h1aa: dout = 8'he0;
    11'h1ab: dout = 8'hfc;
    11'h1ac: dout = 8'h0e;
    11'h1ad: dout = 8'h0e;
    11'h1ae: dout = 8'hfc;
    11'h1af: dout = 8'h00;
    11'h1b0: dout = 8'h7c;
    11'h1b1: dout = 8'he6;
    11'h1b2: dout = 8'he0;
    11'h1b3: dout = 8'hfc;
    11'h1b4: dout = 8'he6;
    11'h1b5: dout = 8'he6;
    11'h1b6: dout = 8'h7c;
    11'h1b7: dout = 8'h00;
    11'h1b8: dout = 8'hfe;
    11'h1b9: dout = 8'h06;
    11'h1ba: dout = 8'h0e;
    11'h1bb: dout = 8'h1c;
    11'h1bc: dout = 8'h38;
    11'h1bd: dout = 8'h38;
    11'h1be: dout = 8'h38;
    11'h1bf: dout = 8'h00;
    11'h1c0: dout = 8'h7c;
    11'h1c1: dout = 8'he6;
    11'h1c2: dout = 8'he6;
    11'h1c3: dout = 8'h7c;
    11'h1c4: dout = 8'he6;
    11'h1c5: dout = 8'he6;
    11'h1c6: dout = 8'h7c;
    11'h1c7: dout = 8'h00;
    11'h1c8: dout = 8'h7c;
    11'h1c9: dout = 8'hce;
    11'h1ca: dout = 8'hce;
    11'h1cb: dout = 8'h7e;
    11'h1cc: dout = 8'h0e;
    11'h1cd: dout = 8'h0e;
    11'h1ce: dout = 8'hfc;
    11'h1cf: dout = 8'h00;
    11'h1d0: dout = 8'h00;
    11'h1d1: dout = 8'h30;
    11'h1d2: dout = 8'h00;
    11'h1d3: dout = 8'h00;
    11'h1d4: dout = 8'h00;
    11'h1d5: dout = 8'h30;
    11'h1d6: dout = 8'h00;
    11'h1d7: dout = 8'h00;
    11'h1d8: dout = 8'h00;
    11'h1d9: dout = 8'h30;
    11'h1da: dout = 8'h00;
    11'h1db: dout = 8'h00;
    11'h1dc: dout = 8'h00;
    11'h1dd: dout = 8'h30;
    11'h1de: dout = 8'h60;
    11'h1df: dout = 8'h00;
    11'h1e0: dout = 8'h00;
    11'h1e1: dout = 8'h18;
    11'h1e2: dout = 8'h30;
    11'h1e3: dout = 8'h60;
    11'h1e4: dout = 8'h30;
    11'h1e5: dout = 8'h18;
    11'h1e6: dout = 8'h00;
    11'h1e7: dout = 8'h00;
    11'h1e8: dout = 8'h00;
    11'h1e9: dout = 8'h00;
    11'h1ea: dout = 8'h7e;
    11'h1eb: dout = 8'h00;
    11'h1ec: dout = 8'h7e;
    11'h1ed: dout = 8'h00;
    11'h1ee: dout = 8'h00;
    11'h1ef: dout = 8'h00;
    11'h1f0: dout = 8'h00;
    11'h1f1: dout = 8'h30;
    11'h1f2: dout = 8'h18;
    11'h1f3: dout = 8'h0c;
    11'h1f4: dout = 8'h18;
    11'h1f5: dout = 8'h30;
    11'h1f6: dout = 8'h00;
    11'h1f7: dout = 8'h00;
    11'h1f8: dout = 8'h7c;
    11'h1f9: dout = 8'hc6;
    11'h1fa: dout = 8'h0e;
    11'h1fb: dout = 8'h1c;
    11'h1fc: dout = 8'h38;
    11'h1fd: dout = 8'h00;
    11'h1fe: dout = 8'h38;
    11'h1ff: dout = 8'h00;
    11'h200: dout = 8'h7c;
    11'h201: dout = 8'hc6;
    11'h202: dout = 8'hde;
    11'h203: dout = 8'hde;
    11'h204: dout = 8'hdc;
    11'h205: dout = 8'hc0;
    11'h206: dout = 8'h7c;
    11'h207: dout = 8'h00;
    11'h208: dout = 8'h7c;
    11'h209: dout = 8'he6;
    11'h20a: dout = 8'he6;
    11'h20b: dout = 8'he6;
    11'h20c: dout = 8'hfe;
    11'h20d: dout = 8'he6;
    11'h20e: dout = 8'he6;
    11'h20f: dout = 8'h00;
    11'h210: dout = 8'hfc;
    11'h211: dout = 8'he6;
    11'h212: dout = 8'he6;
    11'h213: dout = 8'hfc;
    11'h214: dout = 8'he6;
    11'h215: dout = 8'he6;
    11'h216: dout = 8'hfc;
    11'h217: dout = 8'h00;
    11'h218: dout = 8'h7c;
    11'h219: dout = 8'he6;
    11'h21a: dout = 8'he0;
    11'h21b: dout = 8'he0;
    11'h21c: dout = 8'he6;
    11'h21d: dout = 8'he6;
    11'h21e: dout = 8'h7c;
    11'h21f: dout = 8'h00;
    11'h220: dout = 8'hfc;
    11'h221: dout = 8'he6;
    11'h222: dout = 8'he6;
    11'h223: dout = 8'he6;
    11'h224: dout = 8'he6;
    11'h225: dout = 8'he6;
    11'h226: dout = 8'hfc;
    11'h227: dout = 8'h00;
    11'h228: dout = 8'hfe;
    11'h229: dout = 8'he0;
    11'h22a: dout = 8'he0;
    11'h22b: dout = 8'hfe;
    11'h22c: dout = 8'he0;
    11'h22d: dout = 8'he0;
    11'h22e: dout = 8'hfe;
    11'h22f: dout = 8'h00;
    11'h230: dout = 8'hfe;
    11'h231: dout = 8'he0;
    11'h232: dout = 8'he0;
    11'h233: dout = 8'hfe;
    11'h234: dout = 8'he0;
    11'h235: dout = 8'he0;
    11'h236: dout = 8'he0;
    11'h237: dout = 8'h00;
    11'h238: dout = 8'h7c;
    11'h239: dout = 8'he6;
    11'h23a: dout = 8'he0;
    11'h23b: dout = 8'hee;
    11'h23c: dout = 8'he6;
    11'h23d: dout = 8'he6;
    11'h23e: dout = 8'h7c;
    11'h23f: dout = 8'h00;
    11'h240: dout = 8'he6;
    11'h241: dout = 8'he6;
    11'h242: dout = 8'he6;
    11'h243: dout = 8'hfe;
    11'h244: dout = 8'he6;
    11'h245: dout = 8'he6;
    11'h246: dout = 8'he6;
    11'h247: dout = 8'h00;
    11'h248: dout = 8'h38;
    11'h249: dout = 8'h38;
    11'h24a: dout = 8'h38;
    11'h24b: dout = 8'h38;
    11'h24c: dout = 8'h38;
    11'h24d: dout = 8'h38;
    11'h24e: dout = 8'h38;
    11'h24f: dout = 8'h00;
    11'h250: dout = 8'h0e;
    11'h251: dout = 8'h0e;
    11'h252: dout = 8'h0e;
    11'h253: dout = 8'h0e;
    11'h254: dout = 8'hce;
    11'h255: dout = 8'hce;
    11'h256: dout = 8'h7c;
    11'h257: dout = 8'h00;
    11'h258: dout = 8'he6;
    11'h259: dout = 8'hec;
    11'h25a: dout = 8'hf8;
    11'h25b: dout = 8'hf0;
    11'h25c: dout = 8'hf8;
    11'h25d: dout = 8'hec;
    11'h25e: dout = 8'he6;
    11'h25f: dout = 8'h00;
    11'h260: dout = 8'he0;
    11'h261: dout = 8'he0;
    11'h262: dout = 8'he0;
    11'h263: dout = 8'he0;
    11'h264: dout = 8'he0;
    11'h265: dout = 8'he0;
    11'h266: dout = 8'hfe;
    11'h267: dout = 8'h00;
    11'h268: dout = 8'hc6;
    11'h269: dout = 8'hee;
    11'h26a: dout = 8'hfe;
    11'h26b: dout = 8'hd6;
    11'h26c: dout = 8'hc6;
    11'h26d: dout = 8'hc6;
    11'h26e: dout = 8'hc6;
    11'h26f: dout = 8'h00;
    11'h270: dout = 8'hc6;
    11'h271: dout = 8'he6;
    11'h272: dout = 8'hf6;
    11'h273: dout = 8'hfe;
    11'h274: dout = 8'hee;
    11'h275: dout = 8'he6;
    11'h276: dout = 8'he6;
    11'h277: dout = 8'h00;
    11'h278: dout = 8'h7c;
    11'h279: dout = 8'he6;
    11'h27a: dout = 8'he6;
    11'h27b: dout = 8'he6;
    11'h27c: dout = 8'he6;
    11'h27d: dout = 8'he6;
    11'h27e: dout = 8'h7c;
    11'h27f: dout = 8'h00;
    11'h280: dout = 8'hfc;
    11'h281: dout = 8'he6;
    11'h282: dout = 8'he6;
    11'h283: dout = 8'hfc;
    11'h284: dout = 8'he0;
    11'h285: dout = 8'he0;
    11'h286: dout = 8'he0;
    11'h287: dout = 8'h00;
    11'h288: dout = 8'h7c;
    11'h289: dout = 8'he6;
    11'h28a: dout = 8'he6;
    11'h28b: dout = 8'he6;
    11'h28c: dout = 8'he6;
    11'h28d: dout = 8'hea;
    11'h28e: dout = 8'h74;
    11'h28f: dout = 8'h02;
    11'h290: dout = 8'hfc;
    11'h291: dout = 8'he6;
    11'h292: dout = 8'he6;
    11'h293: dout = 8'hfc;
    11'h294: dout = 8'he6;
    11'h295: dout = 8'he6;
    11'h296: dout = 8'he6;
    11'h297: dout = 8'h00;
    11'h298: dout = 8'h7c;
    11'h299: dout = 8'he6;
    11'h29a: dout = 8'he0;
    11'h29b: dout = 8'h7c;
    11'h29c: dout = 8'h0e;
    11'h29d: dout = 8'hce;
    11'h29e: dout = 8'h7c;
    11'h29f: dout = 8'h00;
    11'h2a0: dout = 8'hfe;
    11'h2a1: dout = 8'h38;
    11'h2a2: dout = 8'h38;
    11'h2a3: dout = 8'h38;
    11'h2a4: dout = 8'h38;
    11'h2a5: dout = 8'h38;
    11'h2a6: dout = 8'h38;
    11'h2a7: dout = 8'h00;
    11'h2a8: dout = 8'he6;
    11'h2a9: dout = 8'he6;
    11'h2aa: dout = 8'he6;
    11'h2ab: dout = 8'he6;
    11'h2ac: dout = 8'he6;
    11'h2ad: dout = 8'he6;
    11'h2ae: dout = 8'h7c;
    11'h2af: dout = 8'h00;
    11'h2b0: dout = 8'he6;
    11'h2b1: dout = 8'he6;
    11'h2b2: dout = 8'he6;
    11'h2b3: dout = 8'he6;
    11'h2b4: dout = 8'he6;
    11'h2b5: dout = 8'h7c;
    11'h2b6: dout = 8'h38;
    11'h2b7: dout = 8'h00;
    11'h2b8: dout = 8'hc6;
    11'h2b9: dout = 8'hc6;
    11'h2ba: dout = 8'hc6;
    11'h2bb: dout = 8'hd6;
    11'h2bc: dout = 8'hd6;
    11'h2bd: dout = 8'hfe;
    11'h2be: dout = 8'hfc;
    11'h2bf: dout = 8'h00;
    11'h2c0: dout = 8'he3;
    11'h2c1: dout = 8'h76;
    11'h2c2: dout = 8'h3c;
    11'h2c3: dout = 8'h18;
    11'h2c4: dout = 8'h3c;
    11'h2c5: dout = 8'h6e;
    11'h2c6: dout = 8'hc7;
    11'h2c7: dout = 8'h00;
    11'h2c8: dout = 8'he6;
    11'h2c9: dout = 8'he6;
    11'h2ca: dout = 8'h7c;
    11'h2cb: dout = 8'h38;
    11'h2cc: dout = 8'h38;
    11'h2cd: dout = 8'h38;
    11'h2ce: dout = 8'h38;
    11'h2cf: dout = 8'h00;
    11'h2d0: dout = 8'hfe;
    11'h2d1: dout = 8'h0e;
    11'h2d2: dout = 8'h1c;
    11'h2d3: dout = 8'h38;
    11'h2d4: dout = 8'h70;
    11'h2d5: dout = 8'he0;
    11'h2d6: dout = 8'hfe;
    11'h2d7: dout = 8'h00;
    11'h2d8: dout = 8'h1c;
    11'h2d9: dout = 8'h18;
    11'h2da: dout = 8'h18;
    11'h2db: dout = 8'h18;
    11'h2dc: dout = 8'h18;
    11'h2dd: dout = 8'h18;
    11'h2de: dout = 8'h18;
    11'h2df: dout = 8'h1c;
    11'h2e0: dout = 8'h00;
    11'h2e1: dout = 8'h60;
    11'h2e2: dout = 8'h30;
    11'h2e3: dout = 8'h18;
    11'h2e4: dout = 8'h0c;
    11'h2e5: dout = 8'h06;
    11'h2e6: dout = 8'h03;
    11'h2e7: dout = 8'h00;
    11'h2e8: dout = 8'h70;
    11'h2e9: dout = 8'h30;
    11'h2ea: dout = 8'h30;
    11'h2eb: dout = 8'h30;
    11'h2ec: dout = 8'h30;
    11'h2ed: dout = 8'h30;
    11'h2ee: dout = 8'h30;
    11'h2ef: dout = 8'h70;
    11'h2f0: dout = 8'h18;
    11'h2f1: dout = 8'h3c;
    11'h2f2: dout = 8'h66;
    11'h2f3: dout = 8'hc3;
    11'h2f4: dout = 8'h00;
    11'h2f5: dout = 8'h00;
    11'h2f6: dout = 8'h00;
    11'h2f7: dout = 8'h00;
    11'h2f8: dout = 8'h00;
    11'h2f9: dout = 8'h00;
    11'h2fa: dout = 8'h00;
    11'h2fb: dout = 8'h00;
    11'h2fc: dout = 8'h00;
    11'h2fd: dout = 8'h00;
    11'h2fe: dout = 8'h00;
    11'h2ff: dout = 8'hff;
    11'h300: dout = 8'h30;
    11'h301: dout = 8'h18;
    11'h302: dout = 8'h0c;
    11'h303: dout = 8'h00;
    11'h304: dout = 8'h00;
    11'h305: dout = 8'h00;
    11'h306: dout = 8'h00;
    11'h307: dout = 8'h00;
    11'h308: dout = 8'h00;
    11'h309: dout = 8'h00;
    11'h30a: dout = 8'h7c;
    11'h30b: dout = 8'h0e;
    11'h30c: dout = 8'h7e;
    11'h30d: dout = 8'hce;
    11'h30e: dout = 8'h7e;
    11'h30f: dout = 8'h00;
    11'h310: dout = 8'hc0;
    11'h311: dout = 8'hc0;
    11'h312: dout = 8'hfc;
    11'h313: dout = 8'he6;
    11'h314: dout = 8'he6;
    11'h315: dout = 8'he6;
    11'h316: dout = 8'hfc;
    11'h317: dout = 8'h00;
    11'h318: dout = 8'h00;
    11'h319: dout = 8'h00;
    11'h31a: dout = 8'h7c;
    11'h31b: dout = 8'he6;
    11'h31c: dout = 8'he0;
    11'h31d: dout = 8'he6;
    11'h31e: dout = 8'h7c;
    11'h31f: dout = 8'h00;
    11'h320: dout = 8'h06;
    11'h321: dout = 8'h06;
    11'h322: dout = 8'h7e;
    11'h323: dout = 8'hce;
    11'h324: dout = 8'hce;
    11'h325: dout = 8'hce;
    11'h326: dout = 8'h7e;
    11'h327: dout = 8'h00;
    11'h328: dout = 8'h00;
    11'h329: dout = 8'h00;
    11'h32a: dout = 8'h7c;
    11'h32b: dout = 8'he6;
    11'h32c: dout = 8'hfe;
    11'h32d: dout = 8'he0;
    11'h32e: dout = 8'h7e;
    11'h32f: dout = 8'h00;
    11'h330: dout = 8'h3c;
    11'h331: dout = 8'h70;
    11'h332: dout = 8'h70;
    11'h333: dout = 8'hfc;
    11'h334: dout = 8'h70;
    11'h335: dout = 8'h70;
    11'h336: dout = 8'h70;
    11'h337: dout = 8'h00;
    11'h338: dout = 8'h00;
    11'h339: dout = 8'h00;
    11'h33a: dout = 8'h7c;
    11'h33b: dout = 8'hce;
    11'h33c: dout = 8'hce;
    11'h33d: dout = 8'h7e;
    11'h33e: dout = 8'h0e;
    11'h33f: dout = 8'h7c;
    11'h340: dout = 8'hc0;
    11'h341: dout = 8'hc0;
    11'h342: dout = 8'hfc;
    11'h343: dout = 8'he6;
    11'h344: dout = 8'he6;
    11'h345: dout = 8'he6;
    11'h346: dout = 8'he6;
    11'h347: dout = 8'h00;
    11'h348: dout = 8'h18;
    11'h349: dout = 8'h00;
    11'h34a: dout = 8'h18;
    11'h34b: dout = 8'h38;
    11'h34c: dout = 8'h38;
    11'h34d: dout = 8'h38;
    11'h34e: dout = 8'h38;
    11'h34f: dout = 8'h00;
    11'h350: dout = 8'h0c;
    11'h351: dout = 8'h00;
    11'h352: dout = 8'h0c;
    11'h353: dout = 8'h1c;
    11'h354: dout = 8'h1c;
    11'h355: dout = 8'h1c;
    11'h356: dout = 8'h1c;
    11'h357: dout = 8'hf8;
    11'h358: dout = 8'hc0;
    11'h359: dout = 8'hc0;
    11'h35a: dout = 8'hcc;
    11'h35b: dout = 8'hd8;
    11'h35c: dout = 8'hf0;
    11'h35d: dout = 8'hd8;
    11'h35e: dout = 8'hcc;
    11'h35f: dout = 8'h00;
    11'h360: dout = 8'h18;
    11'h361: dout = 8'h18;
    11'h362: dout = 8'h38;
    11'h363: dout = 8'h38;
    11'h364: dout = 8'h38;
    11'h365: dout = 8'h38;
    11'h366: dout = 8'h38;
    11'h367: dout = 8'h00;
    11'h368: dout = 8'h00;
    11'h369: dout = 8'h00;
    11'h36a: dout = 8'hfc;
    11'h36b: dout = 8'hd6;
    11'h36c: dout = 8'hd6;
    11'h36d: dout = 8'hd6;
    11'h36e: dout = 8'hd6;
    11'h36f: dout = 8'h00;
    11'h370: dout = 8'h00;
    11'h371: dout = 8'h00;
    11'h372: dout = 8'hfc;
    11'h373: dout = 8'he6;
    11'h374: dout = 8'he6;
    11'h375: dout = 8'he6;
    11'h376: dout = 8'he6;
    11'h377: dout = 8'h00;
    11'h378: dout = 8'h00;
    11'h379: dout = 8'h00;
    11'h37a: dout = 8'h7c;
    11'h37b: dout = 8'he6;
    11'h37c: dout = 8'he6;
    11'h37d: dout = 8'he6;
    11'h37e: dout = 8'h7c;
    11'h37f: dout = 8'h00;
    11'h380: dout = 8'h00;
    11'h381: dout = 8'h00;
    11'h382: dout = 8'hfc;
    11'h383: dout = 8'he6;
    11'h384: dout = 8'he6;
    11'h385: dout = 8'hfc;
    11'h386: dout = 8'he0;
    11'h387: dout = 8'he0;
    11'h388: dout = 8'h00;
    11'h389: dout = 8'h00;
    11'h38a: dout = 8'h7e;
    11'h38b: dout = 8'hce;
    11'h38c: dout = 8'hce;
    11'h38d: dout = 8'h7e;
    11'h38e: dout = 8'h0e;
    11'h38f: dout = 8'h0e;
    11'h390: dout = 8'h00;
    11'h391: dout = 8'h00;
    11'h392: dout = 8'hfc;
    11'h393: dout = 8'he6;
    11'h394: dout = 8'he0;
    11'h395: dout = 8'he0;
    11'h396: dout = 8'he0;
    11'h397: dout = 8'h00;
    11'h398: dout = 8'h00;
    11'h399: dout = 8'h00;
    11'h39a: dout = 8'h7e;
    11'h39b: dout = 8'he0;
    11'h39c: dout = 8'h7c;
    11'h39d: dout = 8'h0e;
    11'h39e: dout = 8'hfc;
    11'h39f: dout = 8'h00;
    11'h3a0: dout = 8'h18;
    11'h3a1: dout = 8'h18;
    11'h3a2: dout = 8'h7e;
    11'h3a3: dout = 8'h38;
    11'h3a4: dout = 8'h38;
    11'h3a5: dout = 8'h38;
    11'h3a6: dout = 8'h38;
    11'h3a7: dout = 8'h00;
    11'h3a8: dout = 8'h00;
    11'h3a9: dout = 8'h00;
    11'h3aa: dout = 8'he6;
    11'h3ab: dout = 8'he6;
    11'h3ac: dout = 8'he6;
    11'h3ad: dout = 8'he6;
    11'h3ae: dout = 8'h7e;
    11'h3af: dout = 8'h00;
    11'h3b0: dout = 8'h00;
    11'h3b1: dout = 8'h00;
    11'h3b2: dout = 8'he6;
    11'h3b3: dout = 8'he6;
    11'h3b4: dout = 8'he6;
    11'h3b5: dout = 8'h6c;
    11'h3b6: dout = 8'h38;
    11'h3b7: dout = 8'h00;
    11'h3b8: dout = 8'h00;
    11'h3b9: dout = 8'h00;
    11'h3ba: dout = 8'hd6;
    11'h3bb: dout = 8'hd6;
    11'h3bc: dout = 8'hd6;
    11'h3bd: dout = 8'hd6;
    11'h3be: dout = 8'hfc;
    11'h3bf: dout = 8'h00;
    11'h3c0: dout = 8'h00;
    11'h3c1: dout = 8'h00;
    11'h3c2: dout = 8'he6;
    11'h3c3: dout = 8'h7c;
    11'h3c4: dout = 8'h38;
    11'h3c5: dout = 8'h7c;
    11'h3c6: dout = 8'hce;
    11'h3c7: dout = 8'h00;
    11'h3c8: dout = 8'h00;
    11'h3c9: dout = 8'h00;
    11'h3ca: dout = 8'hce;
    11'h3cb: dout = 8'hce;
    11'h3cc: dout = 8'hce;
    11'h3cd: dout = 8'h7e;
    11'h3ce: dout = 8'h0e;
    11'h3cf: dout = 8'hfc;
    11'h3d0: dout = 8'h00;
    11'h3d1: dout = 8'h00;
    11'h3d2: dout = 8'hfe;
    11'h3d3: dout = 8'h1c;
    11'h3d4: dout = 8'h38;
    11'h3d5: dout = 8'h70;
    11'h3d6: dout = 8'hfe;
    11'h3d7: dout = 8'h00;
    11'h3d8: dout = 8'h0c;
    11'h3d9: dout = 8'h18;
    11'h3da: dout = 8'h18;
    11'h3db: dout = 8'h30;
    11'h3dc: dout = 8'h18;
    11'h3dd: dout = 8'h18;
    11'h3de: dout = 8'h0c;
    11'h3df: dout = 8'h00;
    11'h3e0: dout = 8'h18;
    11'h3e1: dout = 8'h18;
    11'h3e2: dout = 8'h18;
    11'h3e3: dout = 8'h18;
    11'h3e4: dout = 8'h18;
    11'h3e5: dout = 8'h18;
    11'h3e6: dout = 8'h18;
    11'h3e7: dout = 8'h18;
    11'h3e8: dout = 8'h60;
    11'h3e9: dout = 8'h30;
    11'h3ea: dout = 8'h30;
    11'h3eb: dout = 8'h18;
    11'h3ec: dout = 8'h30;
    11'h3ed: dout = 8'h30;
    11'h3ee: dout = 8'h60;
    11'h3ef: dout = 8'h00;
    11'h3f0: dout = 8'h70;
    11'h3f1: dout = 8'hdb;
    11'h3f2: dout = 8'h0e;
    11'h3f3: dout = 8'h00;
    11'h3f4: dout = 8'h00;
    11'h3f5: dout = 8'h00;
    11'h3f6: dout = 8'h00;
    11'h3f7: dout = 8'h00;
    11'h3f8: dout = 8'h00;
    11'h3f9: dout = 8'h00;
    11'h3fa: dout = 8'h10;
    11'h3fb: dout = 8'h28;
    11'h3fc: dout = 8'h44;
    11'h3fd: dout = 8'hfe;
    11'h3fe: dout = 8'h00;
    11'h3ff: dout = 8'h00;
    11'h400: dout = 8'hff;
    11'h401: dout = 8'h80;
    11'h402: dout = 8'h80;
    11'h403: dout = 8'h80;
    11'h404: dout = 8'h80;
    11'h405: dout = 8'h80;
    11'h406: dout = 8'h80;
    11'h407: dout = 8'h80;
    11'h408: dout = 8'hff;
    11'h409: dout = 8'h00;
    11'h40a: dout = 8'h00;
    11'h40b: dout = 8'h00;
    11'h40c: dout = 8'h00;
    11'h40d: dout = 8'h00;
    11'h40e: dout = 8'h00;
    11'h40f: dout = 8'h00;
    11'h410: dout = 8'hff;
    11'h411: dout = 8'h01;
    11'h412: dout = 8'h01;
    11'h413: dout = 8'h01;
    11'h414: dout = 8'h01;
    11'h415: dout = 8'h01;
    11'h416: dout = 8'h01;
    11'h417: dout = 8'h01;
    11'h418: dout = 8'h80;
    11'h419: dout = 8'h80;
    11'h41a: dout = 8'h80;
    11'h41b: dout = 8'h80;
    11'h41c: dout = 8'h80;
    11'h41d: dout = 8'h80;
    11'h41e: dout = 8'h80;
    11'h41f: dout = 8'h80;
    11'h420: dout = 8'h01;
    11'h421: dout = 8'h01;
    11'h422: dout = 8'h01;
    11'h423: dout = 8'h01;
    11'h424: dout = 8'h01;
    11'h425: dout = 8'h01;
    11'h426: dout = 8'h01;
    11'h427: dout = 8'h01;
    11'h428: dout = 8'h80;
    11'h429: dout = 8'h80;
    11'h42a: dout = 8'h80;
    11'h42b: dout = 8'h80;
    11'h42c: dout = 8'h80;
    11'h42d: dout = 8'h80;
    11'h42e: dout = 8'h80;
    11'h42f: dout = 8'hff;
    11'h430: dout = 8'h00;
    11'h431: dout = 8'h00;
    11'h432: dout = 8'h00;
    11'h433: dout = 8'h00;
    11'h434: dout = 8'h00;
    11'h435: dout = 8'h00;
    11'h436: dout = 8'h00;
    11'h437: dout = 8'hff;
    11'h438: dout = 8'h01;
    11'h439: dout = 8'h01;
    11'h43a: dout = 8'h01;
    11'h43b: dout = 8'h01;
    11'h43c: dout = 8'h01;
    11'h43d: dout = 8'h01;
    11'h43e: dout = 8'h01;
    11'h43f: dout = 8'hff;
    11'h440: dout = 8'h80;
    11'h441: dout = 8'h00;
    11'h442: dout = 8'h00;
    11'h443: dout = 8'h00;
    11'h444: dout = 8'h00;
    11'h445: dout = 8'h00;
    11'h446: dout = 8'h00;
    11'h447: dout = 8'h00;
    11'h448: dout = 8'h01;
    11'h449: dout = 8'h00;
    11'h44a: dout = 8'h00;
    11'h44b: dout = 8'h00;
    11'h44c: dout = 8'h00;
    11'h44d: dout = 8'h00;
    11'h44e: dout = 8'h00;
    11'h44f: dout = 8'h00;
    11'h450: dout = 8'h00;
    11'h451: dout = 8'h00;
    11'h452: dout = 8'h00;
    11'h453: dout = 8'h00;
    11'h454: dout = 8'h00;
    11'h455: dout = 8'h00;
    11'h456: dout = 8'h00;
    11'h457: dout = 8'h80;
    11'h458: dout = 8'h00;
    11'h459: dout = 8'h00;
    11'h45a: dout = 8'h00;
    11'h45b: dout = 8'h00;
    11'h45c: dout = 8'h00;
    11'h45d: dout = 8'h00;
    11'h45e: dout = 8'h00;
    11'h45f: dout = 8'h01;
    11'h460: dout = 8'h80;
    11'h461: dout = 8'hc0;
    11'h462: dout = 8'he0;
    11'h463: dout = 8'hf0;
    11'h464: dout = 8'hf8;
    11'h465: dout = 8'hfc;
    11'h466: dout = 8'hfe;
    11'h467: dout = 8'hff;
    11'h468: dout = 8'hff;
    11'h469: dout = 8'h7f;
    11'h46a: dout = 8'h3f;
    11'h46b: dout = 8'h1f;
    11'h46c: dout = 8'h0f;
    11'h46d: dout = 8'h07;
    11'h46e: dout = 8'h03;
    11'h46f: dout = 8'h01;
    11'h470: dout = 8'hff;
    11'h471: dout = 8'hff;
    11'h472: dout = 8'hc0;
    11'h473: dout = 8'hc0;
    11'h474: dout = 8'hc0;
    11'h475: dout = 8'hc0;
    11'h476: dout = 8'hc0;
    11'h477: dout = 8'hc0;
    11'h478: dout = 8'hff;
    11'h479: dout = 8'hff;
    11'h47a: dout = 8'h00;
    11'h47b: dout = 8'h00;
    11'h47c: dout = 8'h00;
    11'h47d: dout = 8'h00;
    11'h47e: dout = 8'h00;
    11'h47f: dout = 8'h00;
    11'h480: dout = 8'hff;
    11'h481: dout = 8'hff;
    11'h482: dout = 8'h03;
    11'h483: dout = 8'h03;
    11'h484: dout = 8'h03;
    11'h485: dout = 8'h03;
    11'h486: dout = 8'h03;
    11'h487: dout = 8'h03;
    11'h488: dout = 8'hc0;
    11'h489: dout = 8'hc0;
    11'h48a: dout = 8'hc0;
    11'h48b: dout = 8'hc0;
    11'h48c: dout = 8'hc0;
    11'h48d: dout = 8'hc0;
    11'h48e: dout = 8'hc0;
    11'h48f: dout = 8'hc0;
    11'h490: dout = 8'h03;
    11'h491: dout = 8'h03;
    11'h492: dout = 8'h03;
    11'h493: dout = 8'h03;
    11'h494: dout = 8'h03;
    11'h495: dout = 8'h03;
    11'h496: dout = 8'h03;
    11'h497: dout = 8'h03;
    11'h498: dout = 8'hc0;
    11'h499: dout = 8'hc0;
    11'h49a: dout = 8'hc0;
    11'h49b: dout = 8'hc0;
    11'h49c: dout = 8'hc0;
    11'h49d: dout = 8'hc0;
    11'h49e: dout = 8'hff;
    11'h49f: dout = 8'hff;
    11'h4a0: dout = 8'h00;
    11'h4a1: dout = 8'h00;
    11'h4a2: dout = 8'h00;
    11'h4a3: dout = 8'h00;
    11'h4a4: dout = 8'h00;
    11'h4a5: dout = 8'h00;
    11'h4a6: dout = 8'hff;
    11'h4a7: dout = 8'hff;
    11'h4a8: dout = 8'h03;
    11'h4a9: dout = 8'h03;
    11'h4aa: dout = 8'h03;
    11'h4ab: dout = 8'h03;
    11'h4ac: dout = 8'h03;
    11'h4ad: dout = 8'h03;
    11'h4ae: dout = 8'hff;
    11'h4af: dout = 8'hff;
    11'h4b0: dout = 8'hc0;
    11'h4b1: dout = 8'hc0;
    11'h4b2: dout = 8'h00;
    11'h4b3: dout = 8'h00;
    11'h4b4: dout = 8'h00;
    11'h4b5: dout = 8'h00;
    11'h4b6: dout = 8'h00;
    11'h4b7: dout = 8'h00;
    11'h4b8: dout = 8'h03;
    11'h4b9: dout = 8'h03;
    11'h4ba: dout = 8'h00;
    11'h4bb: dout = 8'h00;
    11'h4bc: dout = 8'h00;
    11'h4bd: dout = 8'h00;
    11'h4be: dout = 8'h00;
    11'h4bf: dout = 8'h00;
    11'h4c0: dout = 8'h00;
    11'h4c1: dout = 8'h00;
    11'h4c2: dout = 8'h00;
    11'h4c3: dout = 8'h00;
    11'h4c4: dout = 8'h00;
    11'h4c5: dout = 8'h00;
    11'h4c6: dout = 8'hc0;
    11'h4c7: dout = 8'hc0;
    11'h4c8: dout = 8'h00;
    11'h4c9: dout = 8'h00;
    11'h4ca: dout = 8'h00;
    11'h4cb: dout = 8'h00;
    11'h4cc: dout = 8'h00;
    11'h4cd: dout = 8'h00;
    11'h4ce: dout = 8'h03;
    11'h4cf: dout = 8'h03;
    11'h4d0: dout = 8'h00;
    11'h4d1: dout = 8'h00;
    11'h4d2: dout = 8'h00;
    11'h4d3: dout = 8'haa;
    11'h4d4: dout = 8'h00;
    11'h4d5: dout = 8'h00;
    11'h4d6: dout = 8'h00;
    11'h4d7: dout = 8'h00;
    11'h4d8: dout = 8'h00;
    11'h4d9: dout = 8'hfc;
    11'h4da: dout = 8'hfc;
    11'h4db: dout = 8'hfc;
    11'h4dc: dout = 8'hfc;
    11'h4dd: dout = 8'hfc;
    11'h4de: dout = 8'hfc;
    11'h4df: dout = 8'h00;
    11'h4e0: dout = 8'h00;
    11'h4e1: dout = 8'h7e;
    11'h4e2: dout = 8'h7e;
    11'h4e3: dout = 8'h7e;
    11'h4e4: dout = 8'h7e;
    11'h4e5: dout = 8'h7e;
    11'h4e6: dout = 8'h7e;
    11'h4e7: dout = 8'h00;
    11'h4e8: dout = 8'h00;
    11'h4e9: dout = 8'h3f;
    11'h4ea: dout = 8'h3f;
    11'h4eb: dout = 8'h3f;
    11'h4ec: dout = 8'h3f;
    11'h4ed: dout = 8'h3f;
    11'h4ee: dout = 8'h3f;
    11'h4ef: dout = 8'h00;
    11'h4f0: dout = 8'h00;
    11'h4f1: dout = 8'h1f;
    11'h4f2: dout = 8'h1f;
    11'h4f3: dout = 8'h1f;
    11'h4f4: dout = 8'h1f;
    11'h4f5: dout = 8'h1f;
    11'h4f6: dout = 8'h1f;
    11'h4f7: dout = 8'h00;
    11'h4f8: dout = 8'h00;
    11'h4f9: dout = 8'h0f;
    11'h4fa: dout = 8'h0f;
    11'h4fb: dout = 8'h0f;
    11'h4fc: dout = 8'h0f;
    11'h4fd: dout = 8'h0f;
    11'h4fe: dout = 8'h0f;
    11'h4ff: dout = 8'h00;
    11'h500: dout = 8'h00;
    11'h501: dout = 8'h07;
    11'h502: dout = 8'h07;
    11'h503: dout = 8'h07;
    11'h504: dout = 8'h07;
    11'h505: dout = 8'h07;
    11'h506: dout = 8'h07;
    11'h507: dout = 8'h00;
    11'h508: dout = 8'h00;
    11'h509: dout = 8'h03;
    11'h50a: dout = 8'h03;
    11'h50b: dout = 8'h03;
    11'h50c: dout = 8'h03;
    11'h50d: dout = 8'h03;
    11'h50e: dout = 8'h03;
    11'h50f: dout = 8'h00;
    11'h510: dout = 8'h00;
    11'h511: dout = 8'h01;
    11'h512: dout = 8'h01;
    11'h513: dout = 8'h01;
    11'h514: dout = 8'h01;
    11'h515: dout = 8'h01;
    11'h516: dout = 8'h01;
    11'h517: dout = 8'h00;
    11'h518: dout = 8'h00;
    11'h519: dout = 8'h80;
    11'h51a: dout = 8'h80;
    11'h51b: dout = 8'h80;
    11'h51c: dout = 8'h80;
    11'h51d: dout = 8'h80;
    11'h51e: dout = 8'h80;
    11'h51f: dout = 8'h00;
    11'h520: dout = 8'h00;
    11'h521: dout = 8'hc0;
    11'h522: dout = 8'hc0;
    11'h523: dout = 8'hc0;
    11'h524: dout = 8'hc0;
    11'h525: dout = 8'hc0;
    11'h526: dout = 8'hc0;
    11'h527: dout = 8'h00;
    11'h528: dout = 8'h00;
    11'h529: dout = 8'he0;
    11'h52a: dout = 8'he0;
    11'h52b: dout = 8'he0;
    11'h52c: dout = 8'he0;
    11'h52d: dout = 8'he0;
    11'h52e: dout = 8'he0;
    11'h52f: dout = 8'h00;
    11'h530: dout = 8'h00;
    11'h531: dout = 8'hf0;
    11'h532: dout = 8'hf0;
    11'h533: dout = 8'hf0;
    11'h534: dout = 8'hf0;
    11'h535: dout = 8'hf0;
    11'h536: dout = 8'hf0;
    11'h537: dout = 8'h00;
    11'h538: dout = 8'h00;
    11'h539: dout = 8'hf8;
    11'h53a: dout = 8'hf8;
    11'h53b: dout = 8'hf8;
    11'h53c: dout = 8'hf8;
    11'h53d: dout = 8'hf8;
    11'h53e: dout = 8'hf8;
    11'h53f: dout = 8'h00;
    11'h540: dout = 8'haa;
    11'h541: dout = 8'hd6;
    11'h542: dout = 8'haa;
    11'h543: dout = 8'hd6;
    11'h544: dout = 8'haa;
    11'h545: dout = 8'hd6;
    11'h546: dout = 8'haa;
    11'h547: dout = 8'hd6;
    11'h548: dout = 8'hff;
    11'h549: dout = 8'hff;
    11'h54a: dout = 8'h00;
    11'h54b: dout = 8'h00;
    11'h54c: dout = 8'h00;
    11'h54d: dout = 8'h10;
    11'h54e: dout = 8'h38;
    11'h54f: dout = 8'h7c;
    11'h550: dout = 8'hff;
    11'h551: dout = 8'hff;
    11'h552: dout = 8'h00;
    11'h553: dout = 8'h00;
    11'h554: dout = 8'h00;
    11'h555: dout = 8'h00;
    11'h556: dout = 8'h00;
    11'h557: dout = 8'hfe;
    11'h558: dout = 8'hff;
    11'h559: dout = 8'hff;
    11'h55a: dout = 8'h00;
    11'h55b: dout = 8'h00;
    11'h55c: dout = 8'h10;
    11'h55d: dout = 8'h38;
    11'h55e: dout = 8'h7c;
    11'h55f: dout = 8'hfe;
    11'h560: dout = 8'hff;
    11'h561: dout = 8'hff;
    11'h562: dout = 8'h00;
    11'h563: dout = 8'hc3;
    11'h564: dout = 8'he7;
    11'h565: dout = 8'hff;
    11'h566: dout = 8'hdb;
    11'h567: dout = 8'hc3;
    11'h568: dout = 8'h00;
    11'h569: dout = 8'h00;
    11'h56a: dout = 8'h00;
    11'h56b: dout = 8'h00;
    11'h56c: dout = 8'h18;
    11'h56d: dout = 8'h00;
    11'h56e: dout = 8'h00;
    11'h56f: dout = 8'h00;
    11'h570: dout = 8'h00;
    11'h571: dout = 8'hc0;
    11'h572: dout = 8'hc0;
    11'h573: dout = 8'hc0;
    11'h574: dout = 8'hc0;
    11'h575: dout = 8'hc0;
    11'h576: dout = 8'hc0;
    11'h577: dout = 8'hc0;
    11'h578: dout = 8'h00;
    11'h579: dout = 8'hd8;
    11'h57a: dout = 8'hd8;
    11'h57b: dout = 8'hd8;
    11'h57c: dout = 8'hd8;
    11'h57d: dout = 8'hd8;
    11'h57e: dout = 8'hd8;
    11'h57f: dout = 8'hd8;
    11'h580: dout = 8'h00;
    11'h581: dout = 8'hdb;
    11'h582: dout = 8'hdb;
    11'h583: dout = 8'hdb;
    11'h584: dout = 8'hdb;
    11'h585: dout = 8'hdb;
    11'h586: dout = 8'hdb;
    11'h587: dout = 8'hdb;
    11'h588: dout = 8'h00;
    11'h589: dout = 8'h60;
    11'h58a: dout = 8'h60;
    11'h58b: dout = 8'h60;
    11'h58c: dout = 8'h60;
    11'h58d: dout = 8'h60;
    11'h58e: dout = 8'h60;
    11'h58f: dout = 8'h60;
    11'h590: dout = 8'h00;
    11'h591: dout = 8'h6c;
    11'h592: dout = 8'h6c;
    11'h593: dout = 8'h6c;
    11'h594: dout = 8'h6c;
    11'h595: dout = 8'h6c;
    11'h596: dout = 8'h6c;
    11'h597: dout = 8'h6c;
    11'h598: dout = 8'h00;
    11'h599: dout = 8'h6d;
    11'h59a: dout = 8'h6d;
    11'h59b: dout = 8'h6d;
    11'h59c: dout = 8'h6d;
    11'h59d: dout = 8'h6d;
    11'h59e: dout = 8'h6d;
    11'h59f: dout = 8'h6d;
    11'h5a0: dout = 8'h00;
    11'h5a1: dout = 8'h80;
    11'h5a2: dout = 8'h80;
    11'h5a3: dout = 8'h80;
    11'h5a4: dout = 8'h80;
    11'h5a5: dout = 8'h80;
    11'h5a6: dout = 8'h80;
    11'h5a7: dout = 8'h80;
    11'h5a8: dout = 8'h00;
    11'h5a9: dout = 8'hb0;
    11'h5aa: dout = 8'hb0;
    11'h5ab: dout = 8'hb0;
    11'h5ac: dout = 8'hb0;
    11'h5ad: dout = 8'hb0;
    11'h5ae: dout = 8'hb0;
    11'h5af: dout = 8'hb0;
    11'h5b0: dout = 8'h00;
    11'h5b1: dout = 8'hb6;
    11'h5b2: dout = 8'hb6;
    11'h5b3: dout = 8'hb6;
    11'h5b4: dout = 8'hb6;
    11'h5b5: dout = 8'hb6;
    11'h5b6: dout = 8'hb6;
    11'h5b7: dout = 8'hb6;
    11'h5b8: dout = 8'h00;
    11'h5b9: dout = 8'h00;
    11'h5ba: dout = 8'h18;
    11'h5bb: dout = 8'h3c;
    11'h5bc: dout = 8'h3c;
    11'h5bd: dout = 8'h18;
    11'h5be: dout = 8'h00;
    11'h5bf: dout = 8'h00;
    11'h5c0: dout = 8'h00;
    11'h5c1: dout = 8'h00;
    11'h5c2: dout = 8'h00;
    11'h5c3: dout = 8'hf8;
    11'h5c4: dout = 8'h18;
    11'h5c5: dout = 8'hf8;
    11'h5c6: dout = 8'h18;
    11'h5c7: dout = 8'h18;
    11'h5c8: dout = 8'h36;
    11'h5c9: dout = 8'h36;
    11'h5ca: dout = 8'h36;
    11'h5cb: dout = 8'hf6;
    11'h5cc: dout = 8'h06;
    11'h5cd: dout = 8'hf6;
    11'h5ce: dout = 8'h36;
    11'h5cf: dout = 8'h36;
    11'h5d0: dout = 8'h36;
    11'h5d1: dout = 8'h36;
    11'h5d2: dout = 8'h36;
    11'h5d3: dout = 8'h36;
    11'h5d4: dout = 8'h36;
    11'h5d5: dout = 8'h36;
    11'h5d6: dout = 8'h36;
    11'h5d7: dout = 8'h36;
    11'h5d8: dout = 8'h00;
    11'h5d9: dout = 8'h00;
    11'h5da: dout = 8'h00;
    11'h5db: dout = 8'hfe;
    11'h5dc: dout = 8'h06;
    11'h5dd: dout = 8'hf6;
    11'h5de: dout = 8'h36;
    11'h5df: dout = 8'h36;
    11'h5e0: dout = 8'h36;
    11'h5e1: dout = 8'h36;
    11'h5e2: dout = 8'h36;
    11'h5e3: dout = 8'hf6;
    11'h5e4: dout = 8'h06;
    11'h5e5: dout = 8'hfe;
    11'h5e6: dout = 8'h00;
    11'h5e7: dout = 8'h00;
    11'h5e8: dout = 8'h36;
    11'h5e9: dout = 8'h36;
    11'h5ea: dout = 8'h36;
    11'h5eb: dout = 8'hfe;
    11'h5ec: dout = 8'h00;
    11'h5ed: dout = 8'h00;
    11'h5ee: dout = 8'h00;
    11'h5ef: dout = 8'h00;
    11'h5f0: dout = 8'h18;
    11'h5f1: dout = 8'h18;
    11'h5f2: dout = 8'h18;
    11'h5f3: dout = 8'hf8;
    11'h5f4: dout = 8'h18;
    11'h5f5: dout = 8'hf8;
    11'h5f6: dout = 8'h00;
    11'h5f7: dout = 8'h00;
    11'h5f8: dout = 8'h00;
    11'h5f9: dout = 8'h00;
    11'h5fa: dout = 8'h00;
    11'h5fb: dout = 8'hf8;
    11'h5fc: dout = 8'h18;
    11'h5fd: dout = 8'h18;
    11'h5fe: dout = 8'h18;
    11'h5ff: dout = 8'h18;
    11'h600: dout = 8'h18;
    11'h601: dout = 8'h18;
    11'h602: dout = 8'h18;
    11'h603: dout = 8'h1f;
    11'h604: dout = 8'h00;
    11'h605: dout = 8'h00;
    11'h606: dout = 8'h00;
    11'h607: dout = 8'h00;
    11'h608: dout = 8'h18;
    11'h609: dout = 8'h18;
    11'h60a: dout = 8'h18;
    11'h60b: dout = 8'hff;
    11'h60c: dout = 8'h00;
    11'h60d: dout = 8'h00;
    11'h60e: dout = 8'h00;
    11'h60f: dout = 8'h00;
    11'h610: dout = 8'h00;
    11'h611: dout = 8'h00;
    11'h612: dout = 8'h00;
    11'h613: dout = 8'hff;
    11'h614: dout = 8'h18;
    11'h615: dout = 8'h18;
    11'h616: dout = 8'h18;
    11'h617: dout = 8'h18;
    11'h618: dout = 8'h18;
    11'h619: dout = 8'h18;
    11'h61a: dout = 8'h18;
    11'h61b: dout = 8'h1f;
    11'h61c: dout = 8'h18;
    11'h61d: dout = 8'h18;
    11'h61e: dout = 8'h18;
    11'h61f: dout = 8'h18;
    11'h620: dout = 8'h00;
    11'h621: dout = 8'h00;
    11'h622: dout = 8'h00;
    11'h623: dout = 8'hff;
    11'h624: dout = 8'h00;
    11'h625: dout = 8'h00;
    11'h626: dout = 8'h00;
    11'h627: dout = 8'h00;
    11'h628: dout = 8'h18;
    11'h629: dout = 8'h18;
    11'h62a: dout = 8'h18;
    11'h62b: dout = 8'hff;
    11'h62c: dout = 8'h18;
    11'h62d: dout = 8'h18;
    11'h62e: dout = 8'h18;
    11'h62f: dout = 8'h18;
    11'h630: dout = 8'h18;
    11'h631: dout = 8'h18;
    11'h632: dout = 8'h18;
    11'h633: dout = 8'h1f;
    11'h634: dout = 8'h18;
    11'h635: dout = 8'h1f;
    11'h636: dout = 8'h18;
    11'h637: dout = 8'h18;
    11'h638: dout = 8'h36;
    11'h639: dout = 8'h36;
    11'h63a: dout = 8'h36;
    11'h63b: dout = 8'h37;
    11'h63c: dout = 8'h36;
    11'h63d: dout = 8'h36;
    11'h63e: dout = 8'h36;
    11'h63f: dout = 8'h36;
    11'h640: dout = 8'h36;
    11'h641: dout = 8'h36;
    11'h642: dout = 8'h36;
    11'h643: dout = 8'h37;
    11'h644: dout = 8'h30;
    11'h645: dout = 8'h3f;
    11'h646: dout = 8'h00;
    11'h647: dout = 8'h00;
    11'h648: dout = 8'h00;
    11'h649: dout = 8'h00;
    11'h64a: dout = 8'h00;
    11'h64b: dout = 8'h3f;
    11'h64c: dout = 8'h30;
    11'h64d: dout = 8'h37;
    11'h64e: dout = 8'h36;
    11'h64f: dout = 8'h36;
    11'h650: dout = 8'h36;
    11'h651: dout = 8'h36;
    11'h652: dout = 8'h36;
    11'h653: dout = 8'hf7;
    11'h654: dout = 8'h00;
    11'h655: dout = 8'hff;
    11'h656: dout = 8'h00;
    11'h657: dout = 8'h00;
    11'h658: dout = 8'h00;
    11'h659: dout = 8'h00;
    11'h65a: dout = 8'h00;
    11'h65b: dout = 8'hff;
    11'h65c: dout = 8'h00;
    11'h65d: dout = 8'hf7;
    11'h65e: dout = 8'h36;
    11'h65f: dout = 8'h36;
    11'h660: dout = 8'h36;
    11'h661: dout = 8'h36;
    11'h662: dout = 8'h36;
    11'h663: dout = 8'h37;
    11'h664: dout = 8'h30;
    11'h665: dout = 8'h37;
    11'h666: dout = 8'h36;
    11'h667: dout = 8'h36;
    11'h668: dout = 8'h00;
    11'h669: dout = 8'h00;
    11'h66a: dout = 8'h00;
    11'h66b: dout = 8'hff;
    11'h66c: dout = 8'h00;
    11'h66d: dout = 8'hff;
    11'h66e: dout = 8'h00;
    11'h66f: dout = 8'h00;
    11'h670: dout = 8'h36;
    11'h671: dout = 8'h36;
    11'h672: dout = 8'h36;
    11'h673: dout = 8'hf7;
    11'h674: dout = 8'h00;
    11'h675: dout = 8'hf7;
    11'h676: dout = 8'h36;
    11'h677: dout = 8'h36;
    11'h678: dout = 8'h18;
    11'h679: dout = 8'h18;
    11'h67a: dout = 8'h18;
    11'h67b: dout = 8'hff;
    11'h67c: dout = 8'h00;
    11'h67d: dout = 8'hff;
    11'h67e: dout = 8'h00;
    11'h67f: dout = 8'h00;
    11'h680: dout = 8'h36;
    11'h681: dout = 8'h36;
    11'h682: dout = 8'h36;
    11'h683: dout = 8'hff;
    11'h684: dout = 8'h00;
    11'h685: dout = 8'h00;
    11'h686: dout = 8'h00;
    11'h687: dout = 8'h00;
    11'h688: dout = 8'h00;
    11'h689: dout = 8'h00;
    11'h68a: dout = 8'h00;
    11'h68b: dout = 8'hff;
    11'h68c: dout = 8'h00;
    11'h68d: dout = 8'hff;
    11'h68e: dout = 8'h18;
    11'h68f: dout = 8'h18;
    11'h690: dout = 8'h00;
    11'h691: dout = 8'h00;
    11'h692: dout = 8'h00;
    11'h693: dout = 8'hff;
    11'h694: dout = 8'h36;
    11'h695: dout = 8'h36;
    11'h696: dout = 8'h36;
    11'h697: dout = 8'h36;
    11'h698: dout = 8'h36;
    11'h699: dout = 8'h36;
    11'h69a: dout = 8'h36;
    11'h69b: dout = 8'h3f;
    11'h69c: dout = 8'h00;
    11'h69d: dout = 8'h00;
    11'h69e: dout = 8'h00;
    11'h69f: dout = 8'h00;
    11'h6a0: dout = 8'h18;
    11'h6a1: dout = 8'h18;
    11'h6a2: dout = 8'h18;
    11'h6a3: dout = 8'h1f;
    11'h6a4: dout = 8'h18;
    11'h6a5: dout = 8'h1f;
    11'h6a6: dout = 8'h00;
    11'h6a7: dout = 8'h00;
    11'h6a8: dout = 8'h00;
    11'h6a9: dout = 8'h00;
    11'h6aa: dout = 8'h00;
    11'h6ab: dout = 8'h1f;
    11'h6ac: dout = 8'h18;
    11'h6ad: dout = 8'h1f;
    11'h6ae: dout = 8'h18;
    11'h6af: dout = 8'h18;
    11'h6b0: dout = 8'h00;
    11'h6b1: dout = 8'h00;
    11'h6b2: dout = 8'h00;
    11'h6b3: dout = 8'h3f;
    11'h6b4: dout = 8'h36;
    11'h6b5: dout = 8'h36;
    11'h6b6: dout = 8'h36;
    11'h6b7: dout = 8'h36;
    11'h6b8: dout = 8'h36;
    11'h6b9: dout = 8'h36;
    11'h6ba: dout = 8'h36;
    11'h6bb: dout = 8'hff;
    11'h6bc: dout = 8'h36;
    11'h6bd: dout = 8'h36;
    11'h6be: dout = 8'h36;
    11'h6bf: dout = 8'h36;
    11'h6c0: dout = 8'h18;
    11'h6c1: dout = 8'h18;
    11'h6c2: dout = 8'h18;
    11'h6c3: dout = 8'hff;
    11'h6c4: dout = 8'h18;
    11'h6c5: dout = 8'hff;
    11'h6c6: dout = 8'h18;
    11'h6c7: dout = 8'h18;
    11'h6c8: dout = 8'h18;
    11'h6c9: dout = 8'h18;
    11'h6ca: dout = 8'h18;
    11'h6cb: dout = 8'hf8;
    11'h6cc: dout = 8'h00;
    11'h6cd: dout = 8'h00;
    11'h6ce: dout = 8'h00;
    11'h6cf: dout = 8'h00;
    11'h6d0: dout = 8'h00;
    11'h6d1: dout = 8'h00;
    11'h6d2: dout = 8'h00;
    11'h6d3: dout = 8'h1f;
    11'h6d4: dout = 8'h18;
    11'h6d5: dout = 8'h18;
    11'h6d6: dout = 8'h18;
    11'h6d7: dout = 8'h18;
    11'h6d8: dout = 8'hff;
    11'h6d9: dout = 8'hff;
    11'h6da: dout = 8'hff;
    11'h6db: dout = 8'hff;
    11'h6dc: dout = 8'hff;
    11'h6dd: dout = 8'hff;
    11'h6de: dout = 8'hff;
    11'h6df: dout = 8'hff;
    11'h6e0: dout = 8'h00;
    11'h6e1: dout = 8'h00;
    11'h6e2: dout = 8'h00;
    11'h6e3: dout = 8'h00;
    11'h6e4: dout = 8'hff;
    11'h6e5: dout = 8'hff;
    11'h6e6: dout = 8'hff;
    11'h6e7: dout = 8'hff;
    11'h6e8: dout = 8'hf0;
    11'h6e9: dout = 8'hf0;
    11'h6ea: dout = 8'hf0;
    11'h6eb: dout = 8'hf0;
    11'h6ec: dout = 8'hf0;
    11'h6ed: dout = 8'hf0;
    11'h6ee: dout = 8'hf0;
    11'h6ef: dout = 8'hf0;
    11'h6f0: dout = 8'h0f;
    11'h6f1: dout = 8'h0f;
    11'h6f2: dout = 8'h0f;
    11'h6f3: dout = 8'h0f;
    11'h6f4: dout = 8'h0f;
    11'h6f5: dout = 8'h0f;
    11'h6f6: dout = 8'h0f;
    11'h6f7: dout = 8'h0f;
    11'h6f8: dout = 8'hff;
    11'h6f9: dout = 8'hff;
    11'h6fa: dout = 8'hff;
    11'h6fb: dout = 8'hff;
    11'h6fc: dout = 8'h00;
    11'h6fd: dout = 8'h00;
    11'h6fe: dout = 8'h00;
    11'h6ff: dout = 8'h00;
    11'h700: dout = 8'h00;
    11'h701: dout = 8'h00;
    11'h702: dout = 8'h77;
    11'h703: dout = 8'h98;
    11'h704: dout = 8'h98;
    11'h705: dout = 8'h77;
    11'h706: dout = 8'h00;
    11'h707: dout = 8'h00;
    11'h708: dout = 8'h1c;
    11'h709: dout = 8'h36;
    11'h70a: dout = 8'h66;
    11'h70b: dout = 8'hfc;
    11'h70c: dout = 8'hc6;
    11'h70d: dout = 8'hc6;
    11'h70e: dout = 8'hfc;
    11'h70f: dout = 8'hc0;
    11'h710: dout = 8'hfe;
    11'h711: dout = 8'h62;
    11'h712: dout = 8'h60;
    11'h713: dout = 8'h60;
    11'h714: dout = 8'h60;
    11'h715: dout = 8'h60;
    11'h716: dout = 8'h60;
    11'h717: dout = 8'h00;
    11'h718: dout = 8'h00;
    11'h719: dout = 8'h00;
    11'h71a: dout = 8'hff;
    11'h71b: dout = 8'h66;
    11'h71c: dout = 8'h66;
    11'h71d: dout = 8'h66;
    11'h71e: dout = 8'h66;
    11'h71f: dout = 8'h00;
    11'h720: dout = 8'hfe;
    11'h721: dout = 8'h62;
    11'h722: dout = 8'h30;
    11'h723: dout = 8'h18;
    11'h724: dout = 8'h30;
    11'h725: dout = 8'h62;
    11'h726: dout = 8'hfe;
    11'h727: dout = 8'h00;
    11'h728: dout = 8'h00;
    11'h729: dout = 8'h00;
    11'h72a: dout = 8'h3f;
    11'h72b: dout = 8'h66;
    11'h72c: dout = 8'hc6;
    11'h72d: dout = 8'hcc;
    11'h72e: dout = 8'h78;
    11'h72f: dout = 8'h00;
    11'h730: dout = 8'h00;
    11'h731: dout = 8'h00;
    11'h732: dout = 8'h33;
    11'h733: dout = 8'h33;
    11'h734: dout = 8'h33;
    11'h735: dout = 8'h3e;
    11'h736: dout = 8'h30;
    11'h737: dout = 8'hf0;
    11'h738: dout = 8'h00;
    11'h739: dout = 8'h00;
    11'h73a: dout = 8'hff;
    11'h73b: dout = 8'h18;
    11'h73c: dout = 8'h18;
    11'h73d: dout = 8'h18;
    11'h73e: dout = 8'h18;
    11'h73f: dout = 8'h00;
    11'h740: dout = 8'h3c;
    11'h741: dout = 8'h18;
    11'h742: dout = 8'h3c;
    11'h743: dout = 8'h66;
    11'h744: dout = 8'h66;
    11'h745: dout = 8'h3c;
    11'h746: dout = 8'h18;
    11'h747: dout = 8'h3c;
    11'h748: dout = 8'h00;
    11'h749: dout = 8'h7c;
    11'h74a: dout = 8'hc6;
    11'h74b: dout = 8'hfe;
    11'h74c: dout = 8'hc6;
    11'h74d: dout = 8'h7c;
    11'h74e: dout = 8'h00;
    11'h74f: dout = 8'h00;
    11'h750: dout = 8'h00;
    11'h751: dout = 8'h7e;
    11'h752: dout = 8'hc3;
    11'h753: dout = 8'hc3;
    11'h754: dout = 8'hc3;
    11'h755: dout = 8'h66;
    11'h756: dout = 8'he7;
    11'h757: dout = 8'h00;
    11'h758: dout = 8'h1e;
    11'h759: dout = 8'h19;
    11'h75a: dout = 8'h3c;
    11'h75b: dout = 8'h66;
    11'h75c: dout = 8'hc6;
    11'h75d: dout = 8'hcc;
    11'h75e: dout = 8'h78;
    11'h75f: dout = 8'h00;
    11'h760: dout = 8'h00;
    11'h761: dout = 8'h00;
    11'h762: dout = 8'h66;
    11'h763: dout = 8'h99;
    11'h764: dout = 8'h99;
    11'h765: dout = 8'h66;
    11'h766: dout = 8'h00;
    11'h767: dout = 8'h00;
    11'h768: dout = 8'h00;
    11'h769: dout = 8'h03;
    11'h76a: dout = 8'h7c;
    11'h76b: dout = 8'hce;
    11'h76c: dout = 8'he6;
    11'h76d: dout = 8'h7c;
    11'h76e: dout = 8'hc0;
    11'h76f: dout = 8'h00;
    11'h770: dout = 8'h00;
    11'h771: dout = 8'h3e;
    11'h772: dout = 8'hc0;
    11'h773: dout = 8'hfe;
    11'h774: dout = 8'hc0;
    11'h775: dout = 8'h3e;
    11'h776: dout = 8'h00;
    11'h777: dout = 8'h00;
    11'h778: dout = 8'h00;
    11'h779: dout = 8'h7e;
    11'h77a: dout = 8'hc3;
    11'h77b: dout = 8'hc3;
    11'h77c: dout = 8'hc3;
    11'h77d: dout = 8'hc3;
    11'h77e: dout = 8'h00;
    11'h77f: dout = 8'h00;
    11'h780: dout = 8'h00;
    11'h781: dout = 8'hfe;
    11'h782: dout = 8'h00;
    11'h783: dout = 8'hfe;
    11'h784: dout = 8'h00;
    11'h785: dout = 8'hfe;
    11'h786: dout = 8'h00;
    11'h787: dout = 8'h00;
    11'h788: dout = 8'h18;
    11'h789: dout = 8'h18;
    11'h78a: dout = 8'h7e;
    11'h78b: dout = 8'h18;
    11'h78c: dout = 8'h18;
    11'h78d: dout = 8'h7e;
    11'h78e: dout = 8'h00;
    11'h78f: dout = 8'h00;
    11'h790: dout = 8'h70;
    11'h791: dout = 8'h18;
    11'h792: dout = 8'h0c;
    11'h793: dout = 8'h18;
    11'h794: dout = 8'h70;
    11'h795: dout = 8'h00;
    11'h796: dout = 8'hfe;
    11'h797: dout = 8'h00;
    11'h798: dout = 8'h1c;
    11'h799: dout = 8'h30;
    11'h79a: dout = 8'h60;
    11'h79b: dout = 8'h30;
    11'h79c: dout = 8'h1c;
    11'h79d: dout = 8'h00;
    11'h79e: dout = 8'hfe;
    11'h79f: dout = 8'h00;
    11'h7a0: dout = 8'h00;
    11'h7a1: dout = 8'h0e;
    11'h7a2: dout = 8'h1b;
    11'h7a3: dout = 8'h18;
    11'h7a4: dout = 8'h18;
    11'h7a5: dout = 8'h18;
    11'h7a6: dout = 8'h18;
    11'h7a7: dout = 8'h18;
    11'h7a8: dout = 8'h18;
    11'h7a9: dout = 8'h18;
    11'h7aa: dout = 8'h18;
    11'h7ab: dout = 8'h18;
    11'h7ac: dout = 8'h18;
    11'h7ad: dout = 8'hd8;
    11'h7ae: dout = 8'h70;
    11'h7af: dout = 8'h00;
    11'h7b0: dout = 8'h00;
    11'h7b1: dout = 8'h18;
    11'h7b2: dout = 8'h00;
    11'h7b3: dout = 8'h7e;
    11'h7b4: dout = 8'h00;
    11'h7b5: dout = 8'h18;
    11'h7b6: dout = 8'h00;
    11'h7b7: dout = 8'h00;
    11'h7b8: dout = 8'h00;
    11'h7b9: dout = 8'h76;
    11'h7ba: dout = 8'hdc;
    11'h7bb: dout = 8'h00;
    11'h7bc: dout = 8'h76;
    11'h7bd: dout = 8'hdc;
    11'h7be: dout = 8'h00;
    11'h7bf: dout = 8'h00;
    11'h7c0: dout = 8'h3c;
    11'h7c1: dout = 8'h66;
    11'h7c2: dout = 8'h3c;
    11'h7c3: dout = 8'h00;
    11'h7c4: dout = 8'h00;
    11'h7c5: dout = 8'h00;
    11'h7c6: dout = 8'h00;
    11'h7c7: dout = 8'h00;
    11'h7c8: dout = 8'h00;
    11'h7c9: dout = 8'h18;
    11'h7ca: dout = 8'h3c;
    11'h7cb: dout = 8'h18;
    11'h7cc: dout = 8'h00;
    11'h7cd: dout = 8'h00;
    11'h7ce: dout = 8'h00;
    11'h7cf: dout = 8'h00;
    11'h7d0: dout = 8'h00;
    11'h7d1: dout = 8'h00;
    11'h7d2: dout = 8'h00;
    11'h7d3: dout = 8'h00;
    11'h7d4: dout = 8'h18;
    11'h7d5: dout = 8'h00;
    11'h7d6: dout = 8'h00;
    11'h7d7: dout = 8'h00;
    11'h7d8: dout = 8'h0f;
    11'h7d9: dout = 8'h0c;
    11'h7da: dout = 8'h0c;
    11'h7db: dout = 8'h0c;
    11'h7dc: dout = 8'hec;
    11'h7dd: dout = 8'h6c;
    11'h7de: dout = 8'h38;
    11'h7df: dout = 8'h00;
    11'h7e0: dout = 8'hd8;
    11'h7e1: dout = 8'hec;
    11'h7e2: dout = 8'hcc;
    11'h7e3: dout = 8'hcc;
    11'h7e4: dout = 8'h00;
    11'h7e5: dout = 8'h00;
    11'h7e6: dout = 8'h00;
    11'h7e7: dout = 8'h00;
    11'h7e8: dout = 8'hf0;
    11'h7e9: dout = 8'h30;
    11'h7ea: dout = 8'hc0;
    11'h7eb: dout = 8'hf0;
    11'h7ec: dout = 8'h00;
    11'h7ed: dout = 8'h00;
    11'h7ee: dout = 8'h00;
    11'h7ef: dout = 8'h00;
    11'h7f0: dout = 8'h00;
    11'h7f1: dout = 8'h00;
    11'h7f2: dout = 8'h00;
    11'h7f3: dout = 8'h3c;
    11'h7f4: dout = 8'h3c;
    11'h7f5: dout = 8'h3c;
    11'h7f6: dout = 8'h3c;
    11'h7f7: dout = 8'h00;
    11'h7f8: dout = 8'h00;
    11'h7f9: dout = 8'h00;
    11'h7fa: dout = 8'h00;
    11'h7fb: dout = 8'h00;
    11'h7fc: dout = 8'h00;
    11'h7fd: dout = 8'h00;
    11'h7fe: dout = 8'h00;
    11'h7ff: dout = 8'h00;
  endcase
end
endmodule
